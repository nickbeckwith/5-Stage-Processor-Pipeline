`include "cpu.vh"

module cpu(input clk, input rst_n, output hlt, output [15:0] pc_out);
  


endmodule
