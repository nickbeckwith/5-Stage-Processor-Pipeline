module decoder_7_128b(input [6:0] in, output[127:0] out);

  assign out =  (in==7'h00) ? 128'h00000000000000000000000000000001:
                (in==7'h01) ? 128'h00000000000000000000000000000002:
                (in==7'h02) ? 128'h00000000000000000000000000000004:
                (in==7'h03) ? 128'h00000000000000000000000000000008:
                (in==7'h04) ? 128'h00000000000000000000000000000010:
                (in==7'h05) ? 128'h00000000000000000000000000000020:
                (in==7'h06) ? 128'h00000000000000000000000000000040:
                (in==7'h07) ? 128'h00000000000000000000000000000080:
                (in==7'h08) ? 128'h00000000000000000000000000000100:
                (in==7'h09) ? 128'h00000000000000000000000000000200:
                (in==7'h0A) ? 128'h00000000000000000000000000000400:
                (in==7'h0B) ? 128'h00000000000000000000000000000800:
                (in==7'h0C) ? 128'h00000000000000000000000000001000:
                (in==7'h0D) ? 128'h00000000000000000000000000002000:
                (in==7'h0E) ? 128'h00000000000000000000000000004000:
                (in==7'h0F) ? 128'h00000000000000000000000000008000:

                (in==7'h10) ? 128'h00000000000000000000000000010000:
                (in==7'h11) ? 128'h00000000000000000000000000020000:
                (in==7'h12) ? 128'h00000000000000000000000000040000:
                (in==7'h13) ? 128'h00000000000000000000000000080000:
                (in==7'h14) ? 128'h00000000000000000000000000100000:
                (in==7'h15) ? 128'h00000000000000000000000000200000:
                (in==7'h16) ? 128'h00000000000000000000000000400000:
                (in==7'h17) ? 128'h00000000000000000000000000800000:
                (in==7'h18) ? 128'h00000000000000000000000001000000:
                (in==7'h19) ? 128'h00000000000000000000000002000000:
                (in==7'h1A) ? 128'h00000000000000000000000004000000:
                (in==7'h1B) ? 128'h00000000000000000000000008000000:
                (in==7'h1C) ? 128'h00000000000000000000000010000000:
                (in==7'h1D) ? 128'h00000000000000000000000020000000:
                (in==7'h1E) ? 128'h00000000000000000000000040000000:
                (in==7'h1F) ? 128'h00000000000000000000000080000000:

                (in==7'h20) ? 128'h00000000000000000000000100000000:
                (in==7'h21) ? 128'h00000000000000000000000200000000:
                (in==7'h22) ? 128'h00000000000000000000000400000000:
                (in==7'h23) ? 128'h00000000000000000000000800000000:
                (in==7'h24) ? 128'h00000000000000000000001000000000:
                (in==7'h25) ? 128'h00000000000000000000002000000000:
                (in==7'h26) ? 128'h00000000000000000000004000000000:
                (in==7'h27) ? 128'h00000000000000000000008000000000:
                (in==7'h28) ? 128'h00000000000000000000010000000000:
                (in==7'h29) ? 128'h00000000000000000000020000000000:
                (in==7'h2A) ? 128'h00000000000000000000040000000000:
                (in==7'h2B) ? 128'h00000000000000000000080000000000:
                (in==7'h2C) ? 128'h00000000000000000000100000000000:
                (in==7'h2D) ? 128'h00000000000000000000200000000000:
                (in==7'h2E) ? 128'h00000000000000000000400000000000:
                (in==7'h2F) ? 128'h00000000000000000000800000000000:

                (in==7'h30) ? 128'h00000000000000000001000000000000:
                (in==7'h31) ? 128'h00000000000000000002000000000000:
                (in==7'h32) ? 128'h00000000000000000004000000000000:
                (in==7'h33) ? 128'h00000000000000000008000000000000:
                (in==7'h34) ? 128'h00000000000000000010000000000000:
                (in==7'h35) ? 128'h00000000000000000020000000000000:
                (in==7'h36) ? 128'h00000000000000000040000000000000:
                (in==7'h37) ? 128'h00000000000000000080000000000000:
                (in==7'h38) ? 128'h00000000000000000100000000000000:
                (in==7'h39) ? 128'h00000000000000000200000000000000:
                (in==7'h3A) ? 128'h00000000000000000400000000000000:
                (in==7'h3B) ? 128'h00000000000000000800000000000000:
                (in==7'h3C) ? 128'h00000000000000001000000000000000:
                (in==7'h3D) ? 128'h00000000000000002000000000000000:
                (in==7'h3E) ? 128'h00000000000000004000000000000000:
                (in==7'h3F) ? 128'h00000000000000008000000000000000:

                (in==7'h40) ? 128'h00000000000000010000000000000000:
                (in==7'h41) ? 128'h00000000000000020000000000000000:
                (in==7'h42) ? 128'h00000000000000040000000000000000:
                (in==7'h43) ? 128'h00000000000000080000000000000000:
                (in==7'h44) ? 128'h00000000000000100000000000000000:
                (in==7'h45) ? 128'h00000000000000200000000000000000:
                (in==7'h46) ? 128'h00000000000000400000000000000000:
                (in==7'h47) ? 128'h00000000000000800000000000000000:
                (in==7'h48) ? 128'h00000000000001000000000000000000:
                (in==7'h49) ? 128'h00000000000002000000000000000000:
                (in==7'h4A) ? 128'h00000000000004000000000000000000:
                (in==7'h4B) ? 128'h00000000000008000000000000000000:
                (in==7'h4C) ? 128'h00000000000010000000000000000000:
                (in==7'h4D) ? 128'h00000000000020000000000000000000:
                (in==7'h4E) ? 128'h00000000000040000000000000000000:
                (in==7'h4F) ? 128'h00000000000080000000000000000000:

                (in==7'h50) ? 128'h00000000000100000000000000000000:
                (in==7'h51) ? 128'h00000000000200000000000000000000:
                (in==7'h52) ? 128'h00000000000400000000000000000000:
                (in==7'h53) ? 128'h00000000000800000000000000000000:
                (in==7'h54) ? 128'h00000000001000000000000000000000:
                (in==7'h55) ? 128'h00000000002000000000000000000000:
                (in==7'h56) ? 128'h00000000004000000000000000000000:
                (in==7'h57) ? 128'h00000000008000000000000000000000:
                (in==7'h58) ? 128'h00000000010000000000000000000000:
                (in==7'h59) ? 128'h00000000020000000000000000000000:
                (in==7'h5A) ? 128'h00000000040000000000000000000000:
                (in==7'h5B) ? 128'h00000000080000000000000000000000:
                (in==7'h5C) ? 128'h00000000100000000000000000000000:
                (in==7'h5D) ? 128'h00000000200000000000000000000000:
                (in==7'h5E) ? 128'h00000000400000000000000000000000:
                (in==7'h5F) ? 128'h00000000800000000000000000000000:

                (in==7'h60) ? 128'h00000001000000000000000000000000:
                (in==7'h61) ? 128'h00000002000000000000000000000000:
                (in==7'h62) ? 128'h00000004000000000000000000000000:
                (in==7'h63) ? 128'h00000008000000000000000000000000:
                (in==7'h64) ? 128'h00000010000000000000000000000000:
                (in==7'h65) ? 128'h00000020000000000000000000000000:
                (in==7'h66) ? 128'h00000040000000000000000000000000:
                (in==7'h67) ? 128'h00000080000000000000000000000000:
                (in==7'h68) ? 128'h00000100000000000000000000000000:
                (in==7'h69) ? 128'h00000200000000000000000000000000:
                (in==7'h6A) ? 128'h00000400000000000000000000000000:
                (in==7'h6B) ? 128'h00000800000000000000000000000000:
                (in==7'h6C) ? 128'h00001000000000000000000000000000:
                (in==7'h6D) ? 128'h00002000000000000000000000000000:
                (in==7'h6E) ? 128'h00004000000000000000000000000000:
                (in==7'h6F) ? 128'h00008000000000000000000000000000:

                (in==7'h70) ? 128'h00010000000000000000000000000000:
                (in==7'h71) ? 128'h00020000000000000000000000000000:
                (in==7'h72) ? 128'h00040000000000000000000000000000:
                (in==7'h73) ? 128'h00080000000000000000000000000000:
                (in==7'h74) ? 128'h00100000000000000000000000000000:
                (in==7'h75) ? 128'h00200000000000000000000000000000:
                (in==7'h76) ? 128'h00400000000000000000000000000000:
                (in==7'h77) ? 128'h00800000000000000000000000000000:
                (in==7'h78) ? 128'h01000000000000000000000000000000:
                (in==7'h79) ? 128'h02000000000000000000000000000000:
                (in==7'h7A) ? 128'h04000000000000000000000000000000:
                (in==7'h7B) ? 128'h08000000000000000000000000000000:
                (in==7'h7C) ? 128'h10000000000000000000000000000000:
                (in==7'h7D) ? 128'h20000000000000000000000000000000:
                (in==7'h7E) ? 128'h40000000000000000000000000000000:
                (in==7'h7F) ? 128'h80000000000000000000000000000000:
                128'h0;
endmodule
